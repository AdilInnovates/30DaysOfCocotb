// my_module.v
module my_module (
    input wire in_sig,
    output wire out_sig
);
    assign out_sig = in_sig;
endmodule

